/*-------------------------------------------------------------------------------------------
   Digital Direct Synthesizer (DDS)
---------------------------------------------------------------------------------------------
   Author: Fernando Ojeda L.
---------------------------------------------------------------------------------------------
   Description:
---------------------------------------------------------------------------------------------
   DDS that generates a sinewave with 8 bits per sample
   LUT with 256 entries
   
   1. Accumulator with 8-LSB (normal frequency)
   distance between samples = 1 samples
   Period    = (clk*256)
   Frequency = 1/period
   
   
   2. Accumulator with 8-MSB (slower frequency)
   distance between samples = 256 samples (samples are being hold)
   Period    = (clk*256)*256
   Frequency = 1/period
   
---------------------------------------------------------------------------------------------
   Diagram:
---------------------------------------------------------------------------------------------

                   ---> yy - single sinewave
  phase ---> |DDS| ---> y2 - two overlapped sinewaves, low freq + high freq 
                   ---> y3 - impulse response

-------------------------------------------------------------------------------------------*/

module DDS
(
input clk,
input rst,
input  [7:0] phase,
output wire [7:0] yy,
output wire [7:0] y2,
output wire [9:0] y3
);

// *************** Declarations ******************
reg [15:0]  accum;
reg [15:0]  sine;	
reg [15:0]  sine2;	
wire [7:0]  index;
reg  [9:0]  rep;
reg  [9:0]  impulse;


// ************ Accumulator *****************
always@(posedge clk or negedge rst)
begin
	if (rst == 1)
		accum = 16'b0;
	else
		accum = accum + phase;
end

//assign index = accum[15:8]; // take last 8 bits for slower frequency 
assign index  = accum[7:0];   // take first 8 bits for normal frequency


//*****************  Sine LUT ****************************+
always @(posedge clk or negedge rst)
begin
 if (rst == 1) begin
	sine  <= 16'b0;
	sine2 <= 16'b0;
	end
 else begin
 
   // Single Sine LUT
   case (index) 
     8'd  0 : sine <= 16'b               0;  
     8'd  1 : sine <= 16'b      1101000000;  
     8'd  2 : sine <= 16'b     11001000000;  
     8'd  3 : sine <= 16'b    100110000000;  
     8'd  4 : sine <= 16'b    110010000000;  
     8'd  5 : sine <= 16'b    111111000000;  
     8'd  6 : sine <= 16'b   1001011000000;  
     8'd  7 : sine <= 16'b   1010111000000;  
     8'd  8 : sine <= 16'b   1100100000000;  
     8'd  9 : sine <= 16'b   1110000000000;  
     8'd 10 : sine <= 16'b   1111100000000;  
     8'd 11 : sine <= 16'b  10001000000000;  
     8'd 12 : sine <= 16'b  10010100000000;  
     8'd 13 : sine <= 16'b  10100000000000;  
     8'd 14 : sine <= 16'b  10101100000000;  
     8'd 15 : sine <= 16'b  10111000000000;  
     8'd 16 : sine <= 16'b  11000100000000;  
     8'd 17 : sine <= 16'b  11001111000000;  
     8'd 18 : sine <= 16'b  11011011000000;  
     8'd 19 : sine <= 16'b  11100110000000;  
     8'd 20 : sine <= 16'b  11110001000000;  
     8'd 21 : sine <= 16'b  11111100000000;  
     8'd 22 : sine <= 16'b 100000111000000;  
     8'd 23 : sine <= 16'b 100010010000000;  
     8'd 24 : sine <= 16'b 100011100000000;  
     8'd 25 : sine <= 16'b 100100111000000;  
     8'd 26 : sine <= 16'b 100110001000000;  
     8'd 27 : sine <= 16'b 100111011000000;  
     8'd 28 : sine <= 16'b 101000100000000;  
     8'd 29 : sine <= 16'b 101001110000000;  
     8'd 30 : sine <= 16'b 101010111000000;  
     8'd 31 : sine <= 16'b 101100001000000;  
     8'd 32 : sine <= 16'b 101101010000000;  
     8'd 33 : sine <= 16'b 101110010000000;  
     8'd 34 : sine <= 16'b 101111011000000;  
     8'd 35 : sine <= 16'b 110000011000000;  
     8'd 36 : sine <= 16'b 110001011000000;  
     8'd 37 : sine <= 16'b 110010011000000;  
     8'd 38 : sine <= 16'b 110011011000000;  
     8'd 39 : sine <= 16'b 110100010000000;  
     8'd 40 : sine <= 16'b 110101001000000;  
     8'd 41 : sine <= 16'b 110110000000000;  
     8'd 42 : sine <= 16'b 110110111000000;  
     8'd 43 : sine <= 16'b 110111101000000;  
     8'd 44 : sine <= 16'b 111000011000000;  
     8'd 45 : sine <= 16'b 111001001000000;  
     8'd 46 : sine <= 16'b 111001110000000;  
     8'd 47 : sine <= 16'b 111010100000000;  
     8'd 48 : sine <= 16'b 111011001000000;  
     8'd 49 : sine <= 16'b 111011101000000;  
     8'd 50 : sine <= 16'b 111100010000000;  
     8'd 51 : sine <= 16'b 111100110000000;  
     8'd 52 : sine <= 16'b 111101001000000;  
     8'd 53 : sine <= 16'b 111101101000000;  
     8'd 54 : sine <= 16'b 111110000000000;  
     8'd 55 : sine <= 16'b 111110011000000;  
     8'd 56 : sine <= 16'b 111110110000000;  
     8'd 57 : sine <= 16'b 111111000000000;  
     8'd 58 : sine <= 16'b 111111010000000;  
     8'd 59 : sine <= 16'b 111111100000000;  
     8'd 60 : sine <= 16'b 111111101000000;  
     8'd 61 : sine <= 16'b 111111110000000;  
     8'd 62 : sine <= 16'b 111111111000000;  
     8'd 63 : sine <= 16'b 111111111000000;  
     8'd 64 : sine <= 16'b 111111111000000;  
     8'd 65 : sine <= 16'b 111111111000000;  
     8'd 66 : sine <= 16'b 111111111000000;  
     8'd 67 : sine <= 16'b 111111110000000;  
     8'd 68 : sine <= 16'b 111111101000000;  
     8'd 69 : sine <= 16'b 111111100000000;  
     8'd 70 : sine <= 16'b 111111010000000;  
     8'd 71 : sine <= 16'b 111111000000000;  
     8'd 72 : sine <= 16'b 111110110000000;  
     8'd 73 : sine <= 16'b 111110011000000;  
     8'd 74 : sine <= 16'b 111110000000000;  
     8'd 75 : sine <= 16'b 111101101000000;  
     8'd 76 : sine <= 16'b 111101001000000;  
     8'd 77 : sine <= 16'b 111100110000000;  
     8'd 78 : sine <= 16'b 111100010000000;  
     8'd 79 : sine <= 16'b 111011101000000;  
     8'd 80 : sine <= 16'b 111011001000000;  
     8'd 81 : sine <= 16'b 111010100000000;  
     8'd 82 : sine <= 16'b 111001110000000;  
     8'd 83 : sine <= 16'b 111001001000000;  
     8'd 84 : sine <= 16'b 111000011000000;  
     8'd 85 : sine <= 16'b 110111101000000;  
     8'd 86 : sine <= 16'b 110110111000000;  
     8'd 87 : sine <= 16'b 110110000000000;  
     8'd 88 : sine <= 16'b 110101001000000;  
     8'd 89 : sine <= 16'b 110100010000000;  
     8'd 90 : sine <= 16'b 110011011000000;  
     8'd 91 : sine <= 16'b 110010011000000;  
     8'd 92 : sine <= 16'b 110001011000000;  
     8'd 93 : sine <= 16'b 110000011000000;  
     8'd 94 : sine <= 16'b 101111011000000;  
     8'd 95 : sine <= 16'b 101110010000000;  
     8'd 96 : sine <= 16'b 101101010000000;  
     8'd 97 : sine <= 16'b 101100001000000;  
     8'd 98 : sine <= 16'b 101010111000000;  
     8'd 99 : sine <= 16'b 101001110000000;  
     8'd100 : sine <= 16'b 101000100000000;  
     8'd101 : sine <= 16'b 100111011000000;  
     8'd102 : sine <= 16'b 100110001000000;  
     8'd103 : sine <= 16'b 100100111000000;  
     8'd104 : sine <= 16'b 100011100000000;  
     8'd105 : sine <= 16'b 100010010000000;  
     8'd106 : sine <= 16'b 100000111000000;  
     8'd107 : sine <= 16'b  11111100000000;  
     8'd108 : sine <= 16'b  11110001000000;  
     8'd109 : sine <= 16'b  11100110000000;  
     8'd110 : sine <= 16'b  11011011000000;  
     8'd111 : sine <= 16'b  11001111000000;  
     8'd112 : sine <= 16'b  11000100000000;  
     8'd113 : sine <= 16'b  10111000000000;  
     8'd114 : sine <= 16'b  10101100000000;  
     8'd115 : sine <= 16'b  10100000000000;  
     8'd116 : sine <= 16'b  10010100000000;  
     8'd117 : sine <= 16'b  10001000000000;  
     8'd118 : sine <= 16'b   1111100000000;  
     8'd119 : sine <= 16'b   1110000000000;  
     8'd120 : sine <= 16'b   1100100000000;  
     8'd121 : sine <= 16'b   1010111000000;  
     8'd122 : sine <= 16'b   1001011000000;  
     8'd123 : sine <= 16'b    111111000000;  
     8'd124 : sine <= 16'b    110010000000;  
     8'd125 : sine <= 16'b    100110000000;  
     8'd126 : sine <= 16'b     11001000000;  
     8'd127 : sine <= 16'b      1101000000;  
     8'd128 : sine <= 16'b               0;  
     8'd129 : sine <= 16'b1111110011000000;  
     8'd130 : sine <= 16'b1111100111000000;  
     8'd131 : sine <= 16'b1111011010000000;  
     8'd132 : sine <= 16'b1111001110000000;  
     8'd133 : sine <= 16'b1111000001000000;  
     8'd134 : sine <= 16'b1110110101000000;  
     8'd135 : sine <= 16'b1110101001000000;  
     8'd136 : sine <= 16'b1110011100000000;  
     8'd137 : sine <= 16'b1110010000000000;  
     8'd138 : sine <= 16'b1110000100000000;  
     8'd139 : sine <= 16'b1101111000000000;  
     8'd140 : sine <= 16'b1101101100000000;  
     8'd141 : sine <= 16'b1101100000000000;  
     8'd142 : sine <= 16'b1101010100000000;  
     8'd143 : sine <= 16'b1101001000000000;  
     8'd144 : sine <= 16'b1100111100000000;  
     8'd145 : sine <= 16'b1100110001000000;  
     8'd146 : sine <= 16'b1100100101000000;  
     8'd147 : sine <= 16'b1100011010000000;  
     8'd148 : sine <= 16'b1100001111000000;  
     8'd149 : sine <= 16'b1100000100000000;  
     8'd150 : sine <= 16'b1011111001000000;  
     8'd151 : sine <= 16'b1011101110000000;  
     8'd152 : sine <= 16'b1011100100000000;  
     8'd153 : sine <= 16'b1011011001000000;  
     8'd154 : sine <= 16'b1011001111000000;  
     8'd155 : sine <= 16'b1011000101000000;  
     8'd156 : sine <= 16'b1010111100000000;  
     8'd157 : sine <= 16'b1010110010000000;  
     8'd158 : sine <= 16'b1010101001000000;  
     8'd159 : sine <= 16'b1010011111000000;  
     8'd160 : sine <= 16'b1010010110000000;  
     8'd161 : sine <= 16'b1010001110000000;  
     8'd162 : sine <= 16'b1010000101000000;  
     8'd163 : sine <= 16'b1001111101000000;  
     8'd164 : sine <= 16'b1001110101000000;  
     8'd165 : sine <= 16'b1001101101000000;  
     8'd166 : sine <= 16'b1001100101000000;  
     8'd167 : sine <= 16'b1001011110000000;  
     8'd168 : sine <= 16'b1001010111000000;  
     8'd169 : sine <= 16'b1001010000000000;  
     8'd170 : sine <= 16'b1001001001000000;  
     8'd171 : sine <= 16'b1001000011000000;  
     8'd172 : sine <= 16'b1000111101000000;  
     8'd173 : sine <= 16'b1000110111000000;  
     8'd174 : sine <= 16'b1000110010000000;  
     8'd175 : sine <= 16'b1000101100000000;  
     8'd176 : sine <= 16'b1000100111000000;  
     8'd177 : sine <= 16'b1000100011000000;  
     8'd178 : sine <= 16'b1000011110000000;  
     8'd179 : sine <= 16'b1000011010000000;  
     8'd180 : sine <= 16'b1000010111000000;  
     8'd181 : sine <= 16'b1000010011000000;  
     8'd182 : sine <= 16'b1000010000000000;  
     8'd183 : sine <= 16'b1000001101000000;  
     8'd184 : sine <= 16'b1000001010000000;  
     8'd185 : sine <= 16'b1000001000000000;  
     8'd186 : sine <= 16'b1000000110000000;  
     8'd187 : sine <= 16'b1000000100000000;  
     8'd188 : sine <= 16'b1000000011000000;  
     8'd189 : sine <= 16'b1000000010000000;  
     8'd190 : sine <= 16'b1000000001000000;  
     8'd191 : sine <= 16'b1000000001000000;  
     8'd192 : sine <= 16'b1000000001000000;  
     8'd193 : sine <= 16'b1000000001000000;  
     8'd194 : sine <= 16'b1000000001000000;  
     8'd195 : sine <= 16'b1000000010000000;  
     8'd196 : sine <= 16'b1000000011000000;  
     8'd197 : sine <= 16'b1000000100000000;  
     8'd198 : sine <= 16'b1000000110000000;  
     8'd199 : sine <= 16'b1000001000000000;  
     8'd200 : sine <= 16'b1000001010000000;  
     8'd201 : sine <= 16'b1000001101000000;  
     8'd202 : sine <= 16'b1000010000000000;  
     8'd203 : sine <= 16'b1000010011000000;  
     8'd204 : sine <= 16'b1000010111000000;  
     8'd205 : sine <= 16'b1000011010000000;  
     8'd206 : sine <= 16'b1000011110000000;  
     8'd207 : sine <= 16'b1000100011000000;  
     8'd208 : sine <= 16'b1000100111000000;  
     8'd209 : sine <= 16'b1000101100000000;  
     8'd210 : sine <= 16'b1000110010000000;  
     8'd211 : sine <= 16'b1000110111000000;  
     8'd212 : sine <= 16'b1000111101000000;  
     8'd213 : sine <= 16'b1001000011000000;  
     8'd214 : sine <= 16'b1001001001000000;  
     8'd215 : sine <= 16'b1001010000000000;  
     8'd216 : sine <= 16'b1001010111000000;  
     8'd217 : sine <= 16'b1001011110000000;  
     8'd218 : sine <= 16'b1001100101000000;  
     8'd219 : sine <= 16'b1001101101000000;  
     8'd220 : sine <= 16'b1001110101000000;  
     8'd221 : sine <= 16'b1001111101000000;  
     8'd222 : sine <= 16'b1010000101000000;  
     8'd223 : sine <= 16'b1010001110000000;  
     8'd224 : sine <= 16'b1010010110000000;  
     8'd225 : sine <= 16'b1010011111000000;  
     8'd226 : sine <= 16'b1010101001000000;  
     8'd227 : sine <= 16'b1010110010000000;  
     8'd228 : sine <= 16'b1010111100000000;  
     8'd229 : sine <= 16'b1011000101000000;  
     8'd230 : sine <= 16'b1011001111000000;  
     8'd231 : sine <= 16'b1011011001000000;  
     8'd232 : sine <= 16'b1011100100000000;  
     8'd233 : sine <= 16'b1011101110000000;  
     8'd234 : sine <= 16'b1011111001000000;  
     8'd235 : sine <= 16'b1100000100000000;  
     8'd236 : sine <= 16'b1100001111000000;  
     8'd237 : sine <= 16'b1100011010000000;  
     8'd238 : sine <= 16'b1100100101000000;  
     8'd239 : sine <= 16'b1100110001000000;  
     8'd240 : sine <= 16'b1100111100000000;  
     8'd241 : sine <= 16'b1101001000000000;  
     8'd242 : sine <= 16'b1101010100000000;  
     8'd243 : sine <= 16'b1101100000000000;  
     8'd244 : sine <= 16'b1101101100000000;  
     8'd245 : sine <= 16'b1101111000000000;  
     8'd246 : sine <= 16'b1110000100000000;  
     8'd247 : sine <= 16'b1110010000000000;  
     8'd248 : sine <= 16'b1110011100000000;  
     8'd249 : sine <= 16'b1110101001000000;  
     8'd250 : sine <= 16'b1110110101000000;  
     8'd251 : sine <= 16'b1111000001000000;  
     8'd252 : sine <= 16'b1111001110000000;  
     8'd253 : sine <= 16'b1111011010000000;  
     8'd254 : sine <= 16'b1111100111000000;  
     8'd255 : sine <= 16'b1111110011000000;  
   endcase

   // High freq + Low freq Sine LUT
   case (index) 
     8'd  0 : sine2 <= 16'b               0;  
     8'd  1 : sine2 <= 16'b    111101000000;  
     8'd  2 : sine2 <= 16'b     10010000000;  
     8'd  3 : sine2 <= 16'b1111101011000000;  
     8'd  4 : sine2 <= 16'b    101101000000;  
     8'd  5 : sine2 <= 16'b   1100101000000;  
     8'd  6 : sine2 <= 16'b    110101000000;  
     8'd  7 : sine2 <= 16'b     10100000000;  
     8'd  8 : sine2 <= 16'b   1011010000000;  
     8'd  9 : sine2 <= 16'b  10001100000000;  
     8'd 10 : sine2 <= 16'b   1010111000000;  
     8'd 11 : sine2 <= 16'b    111100000000;  
     8'd 12 : sine2 <= 16'b  10000110000000;  
     8'd 13 : sine2 <= 16'b  10110001000000;  
     8'd 14 : sine2 <= 16'b   1111001000000;  
     8'd 15 : sine2 <= 16'b   1100100000000;  
     8'd 16 : sine2 <= 16'b  10110000000000;  
     8'd 17 : sine2 <= 16'b  11010101000000;  
     8'd 18 : sine2 <= 16'b  10011001000000;  
     8'd 19 : sine2 <= 16'b  10001010000000;  
     8'd 20 : sine2 <= 16'b  11011001000000;  
     8'd 21 : sine2 <= 16'b  11110110000000;  
     8'd 22 : sine2 <= 16'b  10111000000000;  
     8'd 23 : sine2 <= 16'b  10110000000000;  
     8'd 24 : sine2 <= 16'b 100000000000000;  
     8'd 25 : sine2 <= 16'b 100010110000000;  
     8'd 26 : sine2 <= 16'b  11010101000000;  
     8'd 27 : sine2 <= 16'b  11010100000000;  
     8'd 28 : sine2 <= 16'b 100100100000000;  
     8'd 29 : sine2 <= 16'b 100110010000000;  
     8'd 30 : sine2 <= 16'b  11110001000000;  
     8'd 31 : sine2 <= 16'b  11110101000000;  
     8'd 32 : sine2 <= 16'b 101000110000000;  
     8'd 33 : sine2 <= 16'b 101001100000000;  
     8'd 34 : sine2 <= 16'b 100001010000000;  
     8'd 35 : sine2 <= 16'b 100010101000000;  
     8'd 36 : sine2 <= 16'b 101100100000000;  
     8'd 37 : sine2 <= 16'b 101100010000000;  
     8'd 38 : sine2 <= 16'b 100100000000000;  
     8'd 39 : sine2 <= 16'b 100110001000000;  
     8'd 40 : sine2 <= 16'b 101111111000000;  
     8'd 41 : sine2 <= 16'b 101110101000000;  
     8'd 42 : sine2 <= 16'b 100110011000000;  
     8'd 43 : sine2 <= 16'b 101001011000000;  
     8'd 44 : sine2 <= 16'b 110010110000000;  
     8'd 45 : sine2 <= 16'b 110000101000000;  
     8'd 46 : sine2 <= 16'b 101000100000000;  
     8'd 47 : sine2 <= 16'b 101100010000000;  
     8'd 48 : sine2 <= 16'b 110101010000000;  
     8'd 49 : sine2 <= 16'b 110010001000000;  
     8'd 50 : sine2 <= 16'b 101010001000000;  
     8'd 51 : sine2 <= 16'b 101110101000000;  
     8'd 52 : sine2 <= 16'b 110111001000000;  
     8'd 53 : sine2 <= 16'b 110011000000000;  
     8'd 54 : sine2 <= 16'b 101011100000000;  
     8'd 55 : sine2 <= 16'b 110000100000000;  
     8'd 56 : sine2 <= 16'b 111000100000000;  
     8'd 57 : sine2 <= 16'b 110011100000000;  
     8'd 58 : sine2 <= 16'b 101100011000000;  
     8'd 59 : sine2 <= 16'b 110010000000000;  
     8'd 60 : sine2 <= 16'b 111001011000000;  
     8'd 61 : sine2 <= 16'b 110011100000000;  
     8'd 62 : sine2 <= 16'b 101100110000000;  
     8'd 63 : sine2 <= 16'b 110011000000000;  
     8'd 64 : sine2 <= 16'b 111001101000000;  
     8'd 65 : sine2 <= 16'b 110011000000000;  
     8'd 66 : sine2 <= 16'b 101100110000000;  
     8'd 67 : sine2 <= 16'b 110011100000000;  
     8'd 68 : sine2 <= 16'b 111001011000000;  
     8'd 69 : sine2 <= 16'b 110010000000000;  
     8'd 70 : sine2 <= 16'b 101100011000000;  
     8'd 71 : sine2 <= 16'b 110011100000000;  
     8'd 72 : sine2 <= 16'b 111000100000000;  
     8'd 73 : sine2 <= 16'b 110000100000000;  
     8'd 74 : sine2 <= 16'b 101011100000000;  
     8'd 75 : sine2 <= 16'b 110011000000000;  
     8'd 76 : sine2 <= 16'b 110111001000000;  
     8'd 77 : sine2 <= 16'b 101110101000000;  
     8'd 78 : sine2 <= 16'b 101010001000000;  
     8'd 79 : sine2 <= 16'b 110010001000000;  
     8'd 80 : sine2 <= 16'b 110101010000000;  
     8'd 81 : sine2 <= 16'b 101100010000000;  
     8'd 82 : sine2 <= 16'b 101000100000000;  
     8'd 83 : sine2 <= 16'b 110000101000000;  
     8'd 84 : sine2 <= 16'b 110010110000000;  
     8'd 85 : sine2 <= 16'b 101001011000000;  
     8'd 86 : sine2 <= 16'b 100110011000000;  
     8'd 87 : sine2 <= 16'b 101110101000000;  
     8'd 88 : sine2 <= 16'b 101111111000000;  
     8'd 89 : sine2 <= 16'b 100110001000000;  
     8'd 90 : sine2 <= 16'b 100100000000000;  
     8'd 91 : sine2 <= 16'b 101100010000000;  
     8'd 92 : sine2 <= 16'b 101100100000000;  
     8'd 93 : sine2 <= 16'b 100010101000000;  
     8'd 94 : sine2 <= 16'b 100001010000000;  
     8'd 95 : sine2 <= 16'b 101001100000000;  
     8'd 96 : sine2 <= 16'b 101000110000000;  
     8'd 97 : sine2 <= 16'b  11110101000000;  
     8'd 98 : sine2 <= 16'b  11110001000000;  
     8'd 99 : sine2 <= 16'b 100110010000000;  
     8'd100 : sine2 <= 16'b 100100100000000;  
     8'd101 : sine2 <= 16'b  11010100000000;  
     8'd102 : sine2 <= 16'b  11010101000000;  
     8'd103 : sine2 <= 16'b 100010110000000;  
     8'd104 : sine2 <= 16'b 100000000000000;  
     8'd105 : sine2 <= 16'b  10110000000000;  
     8'd106 : sine2 <= 16'b  10111000000000;  
     8'd107 : sine2 <= 16'b  11110110000000;  
     8'd108 : sine2 <= 16'b  11011001000000;  
     8'd109 : sine2 <= 16'b  10001010000000;  
     8'd110 : sine2 <= 16'b  10011001000000;  
     8'd111 : sine2 <= 16'b  11010101000000;  
     8'd112 : sine2 <= 16'b  10110000000000;  
     8'd113 : sine2 <= 16'b   1100100000000;  
     8'd114 : sine2 <= 16'b   1111001000000;  
     8'd115 : sine2 <= 16'b  10110001000000;  
     8'd116 : sine2 <= 16'b  10000110000000;  
     8'd117 : sine2 <= 16'b    111100000000;  
     8'd118 : sine2 <= 16'b   1010111000000;  
     8'd119 : sine2 <= 16'b  10001100000000;  
     8'd120 : sine2 <= 16'b   1011010000000;  
     8'd121 : sine2 <= 16'b     10100000000;  
     8'd122 : sine2 <= 16'b    110101000000;  
     8'd123 : sine2 <= 16'b   1100101000000;  
     8'd124 : sine2 <= 16'b    101101000000;  
     8'd125 : sine2 <= 16'b1111101011000000;  
     8'd126 : sine2 <= 16'b     10010000000;  
     8'd127 : sine2 <= 16'b    111101000000;  
     8'd128 : sine2 <= 16'b               0;  
     8'd129 : sine2 <= 16'b1111000011000000;  
     8'd130 : sine2 <= 16'b1111101110000000;  
     8'd131 : sine2 <= 16'b     10101000000;  
     8'd132 : sine2 <= 16'b1111010011000000;  
     8'd133 : sine2 <= 16'b1110011011000000;  
     8'd134 : sine2 <= 16'b1111001011000000;  
     8'd135 : sine2 <= 16'b1111101100000000;  
     8'd136 : sine2 <= 16'b1110100110000000;  
     8'd137 : sine2 <= 16'b1101110100000000;  
     8'd138 : sine2 <= 16'b1110101001000000;  
     8'd139 : sine2 <= 16'b1111000100000000;  
     8'd140 : sine2 <= 16'b1101111010000000;  
     8'd141 : sine2 <= 16'b1101001111000000;  
     8'd142 : sine2 <= 16'b1110000111000000;  
     8'd143 : sine2 <= 16'b1110011100000000;  
     8'd144 : sine2 <= 16'b1101010000000000;  
     8'd145 : sine2 <= 16'b1100101011000000;  
     8'd146 : sine2 <= 16'b1101100111000000;  
     8'd147 : sine2 <= 16'b1101110110000000;  
     8'd148 : sine2 <= 16'b1100100111000000;  
     8'd149 : sine2 <= 16'b1100001010000000;  
     8'd150 : sine2 <= 16'b1101001000000000;  
     8'd151 : sine2 <= 16'b1101010000000000;  
     8'd152 : sine2 <= 16'b1100000000000000;  
     8'd153 : sine2 <= 16'b1011101010000000;  
     8'd154 : sine2 <= 16'b1100101011000000;  
     8'd155 : sine2 <= 16'b1100101100000000;  
     8'd156 : sine2 <= 16'b1011011100000000;  
     8'd157 : sine2 <= 16'b1011001110000000;  
     8'd158 : sine2 <= 16'b1100001111000000;  
     8'd159 : sine2 <= 16'b1100001011000000;  
     8'd160 : sine2 <= 16'b1010111010000000;  
     8'd161 : sine2 <= 16'b1010110100000000;  
     8'd162 : sine2 <= 16'b1011110110000000;  
     8'd163 : sine2 <= 16'b1011101011000000;  
     8'd164 : sine2 <= 16'b1010011100000000;  
     8'd165 : sine2 <= 16'b1010011110000000;  
     8'd166 : sine2 <= 16'b1011100000000000;  
     8'd167 : sine2 <= 16'b1011001111000000;  
     8'd168 : sine2 <= 16'b1010000001000000;  
     8'd169 : sine2 <= 16'b1010001011000000;  
     8'd170 : sine2 <= 16'b1011001101000000;  
     8'd171 : sine2 <= 16'b1010110101000000;  
     8'd172 : sine2 <= 16'b1001101010000000;  
     8'd173 : sine2 <= 16'b1001111011000000;  
     8'd174 : sine2 <= 16'b1010111100000000;  
     8'd175 : sine2 <= 16'b1010011110000000;  
     8'd176 : sine2 <= 16'b1001010110000000;  
     8'd177 : sine2 <= 16'b1001101111000000;  
     8'd178 : sine2 <= 16'b1010101111000000;  
     8'd179 : sine2 <= 16'b1010001011000000;  
     8'd180 : sine2 <= 16'b1001000111000000;  
     8'd181 : sine2 <= 16'b1001101000000000;  
     8'd182 : sine2 <= 16'b1010100100000000;  
     8'd183 : sine2 <= 16'b1001111100000000;  
     8'd184 : sine2 <= 16'b1000111100000000;  
     8'd185 : sine2 <= 16'b1001100100000000;  
     8'd186 : sine2 <= 16'b1010011101000000;  
     8'd187 : sine2 <= 16'b1001110000000000;  
     8'd188 : sine2 <= 16'b1000110101000000;  
     8'd189 : sine2 <= 16'b1001100100000000;  
     8'd190 : sine2 <= 16'b1010011010000000;  
     8'd191 : sine2 <= 16'b1001101000000000;  
     8'd192 : sine2 <= 16'b1000110011000000;  
     8'd193 : sine2 <= 16'b1001101000000000;  
     8'd194 : sine2 <= 16'b1010011010000000;  
     8'd195 : sine2 <= 16'b1001100100000000;  
     8'd196 : sine2 <= 16'b1000110101000000;  
     8'd197 : sine2 <= 16'b1001110000000000;  
     8'd198 : sine2 <= 16'b1010011101000000;  
     8'd199 : sine2 <= 16'b1001100100000000;  
     8'd200 : sine2 <= 16'b1000111100000000;  
     8'd201 : sine2 <= 16'b1001111100000000;  
     8'd202 : sine2 <= 16'b1010100100000000;  
     8'd203 : sine2 <= 16'b1001101000000000;  
     8'd204 : sine2 <= 16'b1001000111000000;  
     8'd205 : sine2 <= 16'b1010001011000000;  
     8'd206 : sine2 <= 16'b1010101111000000;  
     8'd207 : sine2 <= 16'b1001101111000000;  
     8'd208 : sine2 <= 16'b1001010110000000;  
     8'd209 : sine2 <= 16'b1010011110000000;  
     8'd210 : sine2 <= 16'b1010111100000000;  
     8'd211 : sine2 <= 16'b1001111011000000;  
     8'd212 : sine2 <= 16'b1001101010000000;  
     8'd213 : sine2 <= 16'b1010110101000000;  
     8'd214 : sine2 <= 16'b1011001101000000;  
     8'd215 : sine2 <= 16'b1010001011000000;  
     8'd216 : sine2 <= 16'b1010000001000000;  
     8'd217 : sine2 <= 16'b1011001111000000;  
     8'd218 : sine2 <= 16'b1011100000000000;  
     8'd219 : sine2 <= 16'b1010011110000000;  
     8'd220 : sine2 <= 16'b1010011100000000;  
     8'd221 : sine2 <= 16'b1011101011000000;  
     8'd222 : sine2 <= 16'b1011110110000000;  
     8'd223 : sine2 <= 16'b1010110100000000;  
     8'd224 : sine2 <= 16'b1010111010000000;  
     8'd225 : sine2 <= 16'b1100001011000000;  
     8'd226 : sine2 <= 16'b1100001111000000;  
     8'd227 : sine2 <= 16'b1011001110000000;  
     8'd228 : sine2 <= 16'b1011011100000000;  
     8'd229 : sine2 <= 16'b1100101100000000;  
     8'd230 : sine2 <= 16'b1100101011000000;  
     8'd231 : sine2 <= 16'b1011101010000000;  
     8'd232 : sine2 <= 16'b1100000000000000;  
     8'd233 : sine2 <= 16'b1101010000000000;  
     8'd234 : sine2 <= 16'b1101001000000000;  
     8'd235 : sine2 <= 16'b1100001010000000;  
     8'd236 : sine2 <= 16'b1100100111000000;  
     8'd237 : sine2 <= 16'b1101110110000000;  
     8'd238 : sine2 <= 16'b1101100111000000;  
     8'd239 : sine2 <= 16'b1100101011000000;  
     8'd240 : sine2 <= 16'b1101010000000000;  
     8'd241 : sine2 <= 16'b1110011100000000;  
     8'd242 : sine2 <= 16'b1110000111000000;  
     8'd243 : sine2 <= 16'b1101001111000000;  
     8'd244 : sine2 <= 16'b1101111010000000;  
     8'd245 : sine2 <= 16'b1111000100000000;  
     8'd246 : sine2 <= 16'b1110101001000000;  
     8'd247 : sine2 <= 16'b1101110100000000;  
     8'd248 : sine2 <= 16'b1110100110000000;  
     8'd249 : sine2 <= 16'b1111101100000000;  
     8'd250 : sine2 <= 16'b1111001011000000;  
     8'd251 : sine2 <= 16'b1110011011000000;  
     8'd252 : sine2 <= 16'b1111010011000000;  
     8'd253 : sine2 <= 16'b     10101000000;  
     8'd254 : sine2 <= 16'b1111101110000000;  
     8'd255 : sine2 <= 16'b1111000011000000;  
    endcase
  end
end

// **************** impulse response *****************
always@(posedge clk or posedge rst)
begin
if (rst) begin
	   impulse <= 0;
	   rep     <= 0;
	 end
else
	if (rep == 256) begin
	    rep <= 0;
	    impulse <= 10'b0111111111;
	end
	else begin
	    rep <= rep + 1;
	    impulse <= 0;
	end
end


// Outputs
// Scale the sinewaves by 1/256
assign yy = sine[15:8];             // single sinewave
assign y2 = sine2[15:8];            // two overlapped sinewaves, low freq + high freq   
assign y3 = impulse;                // impulse response

endmodule 